* Z:\HOME\ANAGIX\WORK\2020SEPTO\OPAMP\2IN1_TB1.ASC
XX1 NC_01 N003 N004 N003 N006 N001 OUT1 OUT2 2IN1
*V1 N006 0 2.5
*V2 N005 0 SINE(2.5 0.1 1K)
*R1 N001 N005 10K
*R2 N002 N001 100K
*R3 OUT1 N001 100K
*V3 N004 0 5
*V4 N003 0 5

* BLOCK SYMBOL DEFINITIONS 
.SUBCKT 2IN1 VBIAS1 VBIAS2 VDD1 VDD2 VIN+ VIN_ VOUT1 VOUT2
XX1 VIN_ VIN+ VOUT1 VDD1 VBIAS1 0 OPAMP3UREIAUTO
XX2 VIN+ VIN_ VBIAS2 VDD2 VOUT2 0 OPAMP_K_NIIOKA_20200903
.ENDS 2IN1

.SUBCKT OPAMP3UREIAUTO VINM VINP VOUT VDD VBIAS GND
M1 N010 N010 GND GND NMOS L=1U W=16U
M2 N008 N008 N010 GND NMOS L=1U W=16U
M3 N011 N010 GND GND NMOS L=1U W=16U
M4 N007 N008 N011 GND NMOS L=1U W=16U
M5 N001 VBIAS GND GND NMOS L=1U W=34U
M6 N006 VBIAS GND GND NMOS L=1U W=16U
M10 VOUT N009 GND GND NMOS L=1U W=100U
M11 N009 N010 GND GND NMOS L=1U W=16U
M12 VDD N007 N009 GND NMOS L=1U W=16U
M13 N002 N001 VDD VDD PMOS L=1U W=50U
M14 N003 N003 N002 N002 PMOS L=1U W=38U
M15 N006 N006 N003 N003 PMOS L=1U W=38U
M16 N007 N006 N005 N005 PMOS L=1U W=19U
M17 N008 N006 N004 N004 PMOS L=1U W=19U
M18 N004 VINM N002 N002 PMOS L=1U W=25U
M20 VOUT N001 VDD VDD PMOS L=1U W=50U
M21 N005 VINP N002 N002 PMOS L=1U W=25U
M24 N001 N001 VDD VDD PMOS L=1U W=50U
M7 VBIAS VBIAS GND GND NMOS L=1U W=34U
R1 VDD VBIAS 40.25K
C1 VOUT N007 2.9952P
*.INC ./MODELS/OR1_MOS
*.INCLUDE "./BSIM3V3N.MOD"
*.INCLUDE "./BSIM3V3P.MOD"
.ENDS OPAMP3UREIAUTO

.SUBCKT OPAMP_K_NIIOKA_20200903 IN+ IN_ VB VDD OUT GND
M1 N002 N001 VDD VDD PMOS L=3U W=100U
M2 N001 N001 VDD VDD PMOS L=3U W=100U
M4 N001 IN_ N004 GND NMOS L=1U W=400U
M5 N002 IN+ N004 GND NMOS L=1U W=400U
M6 N004 N003 GND GND NMOS L=2.5U W=120U
M7 N003 N003 GND GND NMOS L=2.5U W=10U
M8 OUT N003 GND GND NMOS L=1U W=120U
M3 OUT N002 VDD VDD PMOS L=1U W=240U
C1 N002 OUT 2.9952P
R1 N003 VB 40.25K
*.INCLUDE "./MODELS/OR1_MOS"
.ENDS OPAMP_K_NIIOKA_20200903

.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\ANAGIX\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
.TRAN 10M
.BACKANNO
.END
