* Created by KLayout

* cell 2in1
.SUBCKT 2in1
* net 1 Vin-
* net 2 Vin+
* net 3 Vbia2
* net 4 Vbia1
* net 5 Vout1
* net 6 Vdd1
* net 7 Vdd2
* net 8 Vout2
* net 10 SUBSTRATE
* device instance $1 r0 *1 8.5,72 CAP
C$1 5 9 2.9952e-12
* device instance $2 r0 *1 302,76 CAP
C$2 12 8 2.9952e-12
* device instance $3 r0 *1 170.5,78 HRES
R$3 11 3 40250
* device instance $4 r0 *1 109,141 HRES
R$4 4 6 40250
* device instance $5 r0 *1 154.75,49 NMOS
M$5 10 11 11 10 NMOS L=2.5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $6 r180 *1 271.5,71.5 PMOS
M$6 8 12 7 7 PMOS L=1U W=240U AS=280P AD=280P PS=294U PD=294U
* device instance $12 r0 *1 259,25.5 NMOS
M$12 10 11 8 10 NMOS L=1U W=120U AS=144P AD=144P PS=156U PD=156U
* device instance $17 r180 *1 198.5,79.5 PMOS
M$17 13 13 7 7 PMOS L=3U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $21 m0 *1 220,79.5 PMOS
M$21 12 13 7 7 PMOS L=3U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $25 r180 *1 201,33 NMOS
M$25 13 2 14 10 NMOS L=1U W=400U AS=440P AD=440P PS=462U PD=462U
* device instance $35 r180 *1 241.5,33 NMOS
M$35 12 1 14 10 NMOS L=1U W=400U AS=440P AD=440P PS=462U PD=462U
* device instance $45 r180 *1 159.75,23 NMOS
M$45 14 11 10 10 NMOS L=2.5U W=120U AS=140P AD=140P PS=154U PD=154U
* device instance $51 r0 *1 38.5,61.5 NMOS
M$51 10 15 5 10 NMOS L=1U W=100U AS=200P AD=200P PS=216U PD=216U
* device instance $55 m90 *1 98.5,23 NMOS
M$55 10 4 4 10 NMOS L=1U W=34U AS=68P AD=68P PS=72U PD=72U
* device instance $56 m90 *1 87,23 NMOS
M$56 10 4 20 10 NMOS L=1U W=34U AS=68P AD=68P PS=72U PD=72U
* device instance $57 r0 *1 44.5,30 NMOS
M$57 15 9 6 10 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $58 m90 *1 58,14 NMOS
M$58 10 21 15 10 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $59 m90 *1 65,40.5 NMOS
M$59 24 16 9 10 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $60 r0 *1 72,40.5 NMOS
M$60 21 16 16 10 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $61 r90 *1 95,52 NMOS
M$61 10 4 22 10 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $62 m90 *1 72,14 NMOS
M$62 10 21 21 10 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $63 r0 *1 65,14 NMOS
M$63 10 21 24 10 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $64 r0 *1 60.5,67.5 PMOS
M$64 17 22 9 17 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $65 m90 *1 75,67.5 PMOS
M$65 18 22 16 18 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $66 m90 *1 98.5,104.5 PMOS
M$66 23 19 19 23 PMOS L=1U W=38U AS=76P AD=76P PS=84U PD=84U
* device instance $68 r0 *1 89.5,73.5 PMOS
M$68 19 22 22 19 PMOS L=1U W=38U AS=76P AD=76P PS=84U PD=84U
* device instance $70 r0 *1 62.5,101.5 PMOS
M$70 23 1 17 23 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $71 m90 *1 71.5,101.5 PMOS
M$71 23 2 18 23 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $72 r0 *1 62.5,139 PMOS
M$72 6 20 23 6 PMOS L=1U W=50U AS=100P AD=100P PS=108U PD=108U
* device instance $73 r0 *1 38,139 PMOS
M$73 6 20 5 6 PMOS L=1U W=50U AS=100P AD=100P PS=108U PD=108U
* device instance $74 r0 *1 87.5,139 PMOS
M$74 6 20 20 6 PMOS L=1U W=50U AS=100P AD=100P PS=108U PD=108U
.ENDS 2in1
